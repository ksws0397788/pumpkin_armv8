`include "parameters.h"

module insts_decoder
(
	input [(`INSTS_FETCH_WIDTH_IN_BITS) - 1 : 0]	insts_from_ifetcher_in

);


endmodule
